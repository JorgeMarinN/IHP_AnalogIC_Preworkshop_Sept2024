** sch_path: /home/designer/shared/IHP_AnalogIC_Preworkshop_Sept2024/sg13_cs_amp_full_IHP.sch
**.subckt sg13_cs_amp_full_IHP ref g1 d1 g2 vout
*.ipin ref
*.iopin g1
*.iopin d1
*.iopin g2
*.iopin vout
E1 g1 net1 d1 ref 1000
I0 VDD d1 113.3u
I1 VDD vout 113.3u
XM1 d1 g1 net1 net1 sg13_lv_nmos w=1u l=0.5u ng=1 m=1
XM2 vout g2 net2 net2 sg13_lv_nmos w=1u l=0.5u ng=1 m=1
Vtest2 net2 GND 0
Vtest1 net1 GND 0
**** begin user architecture code

*.option wnflag=1
vds ref 0 0.9
vsup VDD 0 1.8
vin g1 g2 dc=0 ac=60m

cload vout 0 5p

.control
save all

save @n.xm2.nsg13_lv_nmos[gm]
save @n.xm2.nsg13_lv_nmos[ids]
save @n.xm2.nsg13_lv_nmos[gds]

dc vin -0.01 0.01 0.001

let gdsn = @n.xm2.nsg13_lv_nmos[gds]
let gmn = @n.xm2.nsg13_lv_nmos[gm]
let idn = @n.xm2.nsg13_lv_nmos[ids]
let ao = gmn / gdsn

plot deriv(v(vout)) vs v(vout) ao vs v(vout)
plot idn
plot i(vtest1)
plot i(vtest2)
plot v(g2)
plot v(g1)
plot v(d1)

ac dec 100 1 1T
plot vdb(vout)

.endc



.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
