** sch_path: /home/designer/shared/IHP_AnalogIC_Preworkshop_Sept2024/sg13_lv_nmos_charac_IHP.sch
**.subckt sg13_lv_nmos_charac_IHP g1 d1
*.ipin g1
*.iopin d1
XM1 d1 g1 GND GND sg13_lv_nmos w=1.0u l=0.45u ng=5 m=1
**** begin user architecture code



vgs g1 0 dc=0.9
vds d1 0 dc=0.9

.control
save all
*pre_osdi /home/jmarin/Documents/IHP_designs/ihp_design/psp103_nqs.osdi
*  set color0 = white

save @n.xm1.nsg13_lv_nmos[ids]
save @n.xm1.nsg13_lv_nmos[gm]


dc vgs 0 1.8 0.1

let idn = @n.xm1.nsg13_lv_nmos[ids]
let gmn = @n.xm1.nsg13_lv_nmos[gm]
let vthn = @n.xm1.nsg13_lv_nmos[vth]
let vgsn = @n.xm1.nsg13_lv_nmos[vgs]
*let vdsatn = @n.xm1.nsg13_lv_nmos[vdsat]
let vov1 = v(g1) - vthn
let vov2 = 2*idn/gmn

plot idn
plot log(idn)

*let W = 5e-6
*let a = gmn/idn
*setscale a
*plot idn/W
*plot vov2



*wrdata [your_path]/[filename].txt [signals]


.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.GLOBAL GND
.end
